`timescale 1ns / 1ps

    module draw (
      input clk,
      input rst,
      input [9:0] dino_x,
      input [9:0] dino_y,   
      input [9:0] obtacle_x,
      input [9:0] obtacle_y,    
      input [9:0] bird_x,
      input [9:0] bird_y,    
      input [9:0] x,
      input [9:0] y,
      input [1:0]state,
      output reg[11:0]pixel,//12'h0
      output wire dead
    ); 
    parameter dino_w = 10'd40;
    parameter dino_h = 10'd80;
    parameter obtacle_w = 10'd30;
    parameter obtacle_h = 10'd50;
    parameter bird_w = 10'd40;
    parameter bird_h = 10'd30;
     
    wire isobtacle;
    wire isdino;
    wire isbird;
    wire dino_draw;
    wire obtacle_draw;
    wire bird_range;
    wire bird_draw;
    wire black;
    wire sun;
    wire cloud ;
    assign isobtacle = ( x>obtacle_x && x<(obtacle_x+obtacle_w) && y>obtacle_y && y<(obtacle_y+obtacle_h));
    assign isdino = ( x>dino_x && x<(dino_x+dino_w) && y>dino_y && y<(dino_y+dino_h));
    assign isbird = ( x>bird_x && x<(bird_x+bird_w) && y>bird_y && y<(bird_y+bird_h));
    assign dead  = (isobtacle&&isdino&&(state ==2'b01)||isbird&&isdino&&(state ==2'b01));
    assign bird_range = ( x>bird_x && x<(bird_x+bird_w) && y>bird_y && y<(bird_y+10'd2))||
                        ( x>bird_x && x<(bird_x+bird_w) && y>(bird_y+bird_h-10'd2) && y<(bird_y+bird_h))||
                        ( x>bird_x && x<(bird_x+10'd2) && y>bird_y && y<(bird_y+bird_h))||
                        ( x>(bird_x+bird_w-10'd2) && x<(bird_x+bird_w) && y>bird_y && y<(bird_y+bird_h));
    assign cloud =
    ( (x== ( 10'd60)) &&(y > 10'd90) &&(y <10'd100) )||//cloud1
    ( (x== ( 10'd61)) &&(y > 10'd89) &&(y <10'd100) ) ||
    ( (x== ( 10'd62)) &&(y > 10'd90) &&(y <10'd100) )||
    ( (x== ( 10'd63)) &&(y > 10'd87) &&(y <10'd100) ) ||
    ( (x== ( 10'd64)) &&(y > 10'd86) &&(y <10'd100) )||
    ( (x== ( 10'd65)) &&(y > 10'd87) &&(y <10'd100) ) ||
    ( (x== ( 10'd66)) &&(y > 10'd84) &&(y <10'd100) )||
    ( (x== ( 10'd67)) &&(y > 10'd83) &&(y <10'd100) ) ||
    ( (x== ( 10'd68)) &&(y > 10'd84) &&(y <10'd100) )||
    ( (x== ( 10'd69)) &&(y > 10'd82) &&(y <10'd100) ) ||
    ( (x== ( 10'd70)) &&(y > 10'd81) &&(y <10'd100) )||
    ( (x== ( 10'd71)) &&(y > 10'd82) &&(y <10'd100) ) ||
    ( (x== ( 10'd72)) &&(y > 10'd79) &&(y <10'd100) )||
    ( (x== ( 10'd73)) &&(y > 10'd78) &&(y <10'd100) ) ||
    ( (x== ( 10'd74)) &&(y > 10'd79) &&(y <10'd100) )||
    ( (x== ( 10'd75)) &&(y > 10'd78) &&(y <10'd100) ) ||
    ( (x== ( 10'd76)) &&(y > 10'd77) &&(y <10'd100) )||
    ( (x== ( 10'd77)) &&(y > 10'd78) &&(y <10'd100) ) ||
    ( (x== ( 10'd78)) &&(y > 10'd81) &&(y <10'd100) )||
    ( (x== ( 10'd79)) &&(y > 10'd80) &&(y <10'd100) ) ||
    ( (x== ( 10'd80)) &&(y > 10'd81) &&(y <10'd100) )||
    ( (x== ( 10'd81)) &&(y > 10'd82) &&(y <10'd100) ) ||
    ( (x== ( 10'd82)) &&(y > 10'd81) &&(y <10'd100) )||
    ( (x== ( 10'd83)) &&(y > 10'd82) &&(y <10'd100) ) ||
    ( (x== ( 10'd84)) &&(y > 10'd82) &&(y <10'd100) )||
    ( (x== ( 10'd85)) &&(y > 10'd85) &&(y <10'd100) ) ||
    ( (x== ( 10'd86)) &&(y > 10'd84) &&(y <10'd100) )||
    ( (x== ( 10'd87)) &&(y > 10'd85) &&(y <10'd100) ) ||
    ( (x== ( 10'd88)) &&(y > 10'd83) &&(y <10'd100) )||
    ( (x== ( 10'd89)) &&(y > 10'd83) &&(y <10'd100) ) ||
    ( (x== ( 10'd90)) &&(y > 10'd82) &&(y <10'd100) )||
    ( (x== ( 10'd91)) &&(y > 10'd83) &&(y <10'd100) ) ||
    ( (x== ( 10'd92)) &&(y > 10'd85) &&(y <10'd100) )||
    ( (x== ( 10'd93)) &&(y > 10'd84) &&(y <10'd100) ) ||
    ( (x== ( 10'd94)) &&(y > 10'd85) &&(y <10'd100) )||
    ( (x== ( 10'd95)) &&(y > 10'd86) &&(y <10'd100) ) ||
    ( (x== ( 10'd96)) &&(y > 10'd85) &&(y <10'd100) )||
    ( (x== ( 10'd97)) &&(y > 10'd86) &&(y <10'd100) ) ||
    ( (x== ( 10'd98)) &&(y > 10'd88) &&(y <10'd100) )||
    ( (x== ( 10'd99)) &&(y > 10'd87) &&(y <10'd100) ) ||
    ( (x== ( 10'd100)) &&(y > 10'd88) &&(y <10'd100) )||
    ( (x== ( 10'd101)) &&(y > 10'd87) &&(y <10'd100) ) ||
    ( (x== ( 10'd102)) &&(y > 10'd86) &&(y <10'd100) )||
    ( (x== ( 10'd103)) &&(y > 10'd87) &&(y <10'd100) ) ||
    ( (x== ( 10'd104)) &&(y > 10'd88) &&(y <10'd100) )||
    ( (x== ( 10'd105)) &&(y > 10'd87) &&(y <10'd100) ) ||
    ( (x== ( 10'd106)) &&(y > 10'd88) &&(y <10'd100) )||
    ( (x== ( 10'd107)) &&(y > 10'd86) &&(y <10'd100) ) ||
    ( (x== ( 10'd108)) &&(y > 10'd85) &&(y <10'd100) )||
    ( (x== ( 10'd109)) &&(y > 10'd85) &&(y <10'd100) ) ||
    ( (x== ( 10'd110)) &&(y > 10'd86) &&(y <10'd100) )||
    ( (x== ( 10'd111)) &&(y > 10'd83) &&(y <10'd100) ) ||
    ( (x== ( 10'd112)) &&(y > 10'd82) &&(y <10'd100) )||
    ( (x== ( 10'd113)) &&(y > 10'd83) &&(y <10'd100) ) ||
    ( (x== ( 10'd114)) &&(y > 10'd81) &&(y <10'd100) )||
    ( (x== ( 10'd115)) &&(y > 10'd80) &&(y <10'd100) ) ||
    ( (x== ( 10'd116)) &&(y > 10'd81) &&(y <10'd100) )||
    ( (x== ( 10'd117)) &&(y > 10'd79) &&(y <10'd100) ) ||
    ( (x== ( 10'd118)) &&(y > 10'd78) &&(y <10'd100) )||
    ( (x== ( 10'd119)) &&(y > 10'd79) &&(y <10'd100) ) ||
    ( (x== ( 10'd120)) &&(y > 10'd79) &&(y <10'd100) ) ||
    ( (y== ( 10'd91)) &&(x > 10'd57) &&(x <10'd60) ) ||//cloud1_left
    ( (y== ( 10'd92)) &&(x > 10'd56) &&(x <10'd60) ) ||
    ( (y== ( 10'd93)) &&(x > 10'd57) &&(x <10'd60) ) ||
    ( (y== ( 10'd94)) &&(x > 10'd56) &&(x <10'd60) ) ||
    ( (y== ( 10'd95)) &&(x > 10'd57) &&(x <10'd60) ) ||
    ( (y== ( 10'd96)) &&(x > 10'd56) &&(x <10'd60) ) ||
    ( (y== ( 10'd97)) &&(x > 10'd54) &&(x <10'd60) ) ||
    ( (y== ( 10'd98)) &&(x > 10'd55) &&(x <10'd60) ) ||
    ( (y== ( 10'd99)) &&(x > 10'd54) &&(x <10'd60) ) ||
    ( (y== ( 10'd80)) &&(x > 10'd120) &&(x <10'd122) ) ||//cloud1_right
    ( (y== ( 10'd81)) &&(x > 10'd120) &&(x <10'd121) ) ||
    ( (y== ( 10'd82)) &&(x > 10'd120) &&(x <10'd122) ) ||
    ( (y== ( 10'd83)) &&(x > 10'd120) &&(x <10'd123) ) ||
    ( (y== ( 10'd84)) &&(x > 10'd120) &&(x <10'd122) ) ||
    ( (y== ( 10'd85)) &&(x > 10'd120) &&(x <10'd123) ) ||
    ( (y== ( 10'd86)) &&(x > 10'd120) &&(x <10'd123) ) ||
    ( (y== ( 10'd87)) &&(x > 10'd120) &&(x <10'd124) ) ||
    ( (y== ( 10'd88)) &&(x > 10'd120) &&(x <10'd123) ) ||
    ( (y== ( 10'd89)) &&(x > 10'd120) &&(x <10'd124) ) ||
    ( (y== ( 10'd90)) &&(x > 10'd120) &&(x <10'd123) ) ||
    ( (y== ( 10'd91)) &&(x > 10'd120) &&(x <10'd123) ) ||
    ( (y== ( 10'd92)) &&(x > 10'd120) &&(x <10'd122) ) ||
    ( (y== ( 10'd93)) &&(x > 10'd120) &&(x <10'd123) ) ||
    ( (y== ( 10'd94)) &&(x > 10'd120) &&(x <10'd125) ) ||
    ( (y== ( 10'd95)) &&(x > 10'd120) &&(x <10'd124) ) ||
    ( (y== ( 10'd96)) &&(x > 10'd120) &&(x <10'd125) ) ||
    ( (y== ( 10'd97)) &&(x > 10'd120) &&(x <10'd126) ) ||
    ( (y== ( 10'd98)) &&(x > 10'd120) &&(x <10'd125) ) ||
    ( (y== ( 10'd99)) &&(x > 10'd120) &&(x <10'd126) ) ||
    ( (x== ( 10'd130)) &&(y > 10'd160) &&(y <10'd170) )||//cloud2
    ( (x== ( 10'd131)) &&(y > 10'd157) &&(y <10'd170) ) ||
    ( (x== ( 10'd132)) &&(y > 10'd160) &&(y <10'd170) )||
    ( (x== ( 10'd133)) &&(y > 10'd157) &&(y <10'd170) ) ||
    ( (x== ( 10'd134)) &&(y > 10'd156) &&(y <10'd170) )||
    ( (x== ( 10'd135)) &&(y > 10'd157) &&(y <10'd170) ) ||
    ( (x== ( 10'd136)) &&(y > 10'd154) &&(y <10'd170) )||
    ( (x== ( 10'd137)) &&(y > 10'd153) &&(y <10'd170) ) ||
    ( (x== ( 10'd138)) &&(y > 10'd154) &&(y <10'd170) )||
    ( (x== ( 10'd139)) &&(y > 10'd152) &&(y <10'd170) ) ||
    ( (x== ( 10'd140)) &&(y > 10'd151) &&(y <10'd170) )||
    ( (x== ( 10'd141)) &&(y > 10'd152) &&(y <10'd170) ) ||
    ( (x== ( 10'd142)) &&(y > 10'd149) &&(y <10'd170) )||
    ( (x== ( 10'd143)) &&(y > 10'd148) &&(y <10'd170) ) ||
    ( (x== ( 10'd144)) &&(y > 10'd149) &&(y <10'd170) )||
    ( (x== ( 10'd145)) &&(y > 10'd148) &&(y <10'd170) ) ||
    ( (x== ( 10'd146)) &&(y > 10'd147) &&(y <10'd170) )||
    ( (x== ( 10'd147)) &&(y > 10'd148) &&(y <10'd170) ) ||
    ( (x== ( 10'd148)) &&(y > 10'd151) &&(y <10'd170) )||
    ( (x== ( 10'd149)) &&(y > 10'd150) &&(y <10'd170) ) ||
    ( (x== ( 10'd150)) &&(y > 10'd151) &&(y <10'd170) )||
    ( (x== ( 10'd151)) &&(y > 10'd152) &&(y <10'd170) ) ||
    ( (x== ( 10'd152)) &&(y > 10'd151) &&(y <10'd170) )||
    ( (x== ( 10'd153)) &&(y > 10'd152) &&(y <10'd170) ) ||
    ( (x== ( 10'd154)) &&(y > 10'd152) &&(y <10'd170) )||
    ( (x== ( 10'd155)) &&(y > 10'd155) &&(y <10'd170) ) ||
    ( (x== ( 10'd156)) &&(y > 10'd154) &&(y <10'd170) )||
    ( (x== ( 10'd157)) &&(y > 10'd155) &&(y <10'd170) ) ||
    ( (x== ( 10'd158)) &&(y > 10'd153) &&(y <10'd170) )||
    ( (x== ( 10'd159)) &&(y > 10'd153) &&(y <10'd170) ) ||
    ( (x== ( 10'd160)) &&(y > 10'd152) &&(y <10'd170) )||
    ( (x== ( 10'd161)) &&(y > 10'd153) &&(y <10'd170) ) ||
    ( (x== ( 10'd162)) &&(y > 10'd155) &&(y <10'd170) )||
    ( (x== ( 10'd163)) &&(y > 10'd154) &&(y <10'd170) ) ||
    ( (x== ( 10'd164)) &&(y > 10'd155) &&(y <10'd170) )||
    ( (x== ( 10'd165)) &&(y > 10'd156) &&(y <10'd170) ) ||
    ( (x== ( 10'd166)) &&(y > 10'd155) &&(y <10'd170) )||
    ( (x== ( 10'd167)) &&(y > 10'd156) &&(y <10'd170) ) ||
    ( (x== ( 10'd168)) &&(y > 10'd158) &&(y <10'd170) )||
    ( (x== ( 10'd169)) &&(y > 10'd157) &&(y <10'd170) ) ||
    ( (x== ( 10'd170)) &&(y > 10'd158) &&(y <10'd170) )||
    ( (x== ( 10'd171)) &&(y > 10'd157) &&(y <10'd170) ) ||
    ( (x== ( 10'd172)) &&(y > 10'd156) &&(y <10'd170) )||
    ( (x== ( 10'd173)) &&(y > 10'd157) &&(y <10'd170) ) ||
    ( (x== ( 10'd174)) &&(y > 10'd158) &&(y <10'd170) )||
    ( (x== ( 10'd175)) &&(y > 10'd157) &&(y <10'd170) ) ||
    ( (x== ( 10'd176)) &&(y > 10'd158) &&(y <10'd170) )||
    ( (x== ( 10'd177)) &&(y > 10'd156) &&(y <10'd170) ) ||
    ( (x== ( 10'd178)) &&(y > 10'd155) &&(y <10'd170) )||
    ( (x== ( 10'd179)) &&(y > 10'd155) &&(y <10'd170) ) ||
    ( (x== ( 10'd180)) &&(y > 10'd156) &&(y <10'd170) )||
    ( (x== ( 10'd181)) &&(y > 10'd153) &&(y <10'd170) ) ||
    ( (x== ( 10'd182)) &&(y > 10'd152) &&(y <10'd170) )||
    ( (x== ( 10'd183)) &&(y > 10'd153) &&(y <10'd170) ) ||
    ( (x== ( 10'd184)) &&(y > 10'd151) &&(y <10'd170) )||
    ( (x== ( 10'd185)) &&(y > 10'd150) &&(y <10'd170) ) ||
    ( (x== ( 10'd186)) &&(y > 10'd151) &&(y <10'd170) )||
    ( (x== ( 10'd187)) &&(y > 10'd149) &&(y <10'd170) ) ||
    ( (x== ( 10'd188)) &&(y > 10'd148) &&(y <10'd170) )||
    ( (x== ( 10'd189)) &&(y > 10'd149) &&(y <10'd170) ) ||
    ( (x== ( 10'd190)) &&(y > 10'd149) &&(y <10'd100) ) ||
    ( (y== ( 10'd161)) &&(x > 10'd127) &&(x <10'd130) ) ||//cloud2_left
    ( (y== ( 10'd162)) &&(x > 10'd126) &&(x <10'd130) ) ||
    ( (y== ( 10'd163)) &&(x > 10'd127) &&(x <10'd130) ) ||
    ( (y== ( 10'd164)) &&(x > 10'd126) &&(x <10'd130) ) ||
    ( (y== ( 10'd165)) &&(x > 10'd127) &&(x <10'd130) ) ||
    ( (y== ( 10'd166)) &&(x > 10'd126) &&(x <10'd130) ) ||
    ( (y== ( 10'd167)) &&(x > 10'd124) &&(x <10'd130) ) ||
    ( (y== ( 10'd168)) &&(x > 10'd125) &&(x <10'd130) ) ||
    ( (y== ( 10'd169)) &&(x > 10'd124) &&(x <10'd130) ) ||
    ( (y== ( 10'd150)) &&(x > 10'd189) &&(x <10'd192) ) ||//cloud2_right
    ( (y== ( 10'd151)) &&(x > 10'd189) &&(x <10'd191) ) ||
    ( (y== ( 10'd152)) &&(x > 10'd189) &&(x <10'd192) ) ||
    ( (y== ( 10'd153)) &&(x > 10'd189) &&(x <10'd193) ) ||
    ( (y== ( 10'd154)) &&(x > 10'd189) &&(x <10'd192) ) ||
    ( (y== ( 10'd155)) &&(x > 10'd189) &&(x <10'd193) ) ||
    ( (y== ( 10'd156)) &&(x > 10'd189) &&(x <10'd193) ) ||
    ( (y== ( 10'd157)) &&(x > 10'd189) &&(x <10'd194) ) ||
    ( (y== ( 10'd158)) &&(x > 10'd189) &&(x <10'd193) ) ||
    ( (y== ( 10'd159)) &&(x > 10'd189) &&(x <10'd194) ) ||
    ( (y== ( 10'd160)) &&(x > 10'd189) &&(x <10'd193) ) ||
    ( (y== ( 10'd161)) &&(x > 10'd189) &&(x <10'd193) ) ||
    ( (y== ( 10'd162)) &&(x > 10'd189) &&(x <10'd192) ) ||
    ( (y== ( 10'd163)) &&(x > 10'd189) &&(x <10'd193) ) ||
    ( (y== ( 10'd164)) &&(x > 10'd189) &&(x <10'd195) ) ||
    ( (y== ( 10'd165)) &&(x > 10'd189) &&(x <10'd194) ) ||
    ( (y== ( 10'd166)) &&(x > 10'd189) &&(x <10'd195) ) ||
    ( (y== ( 10'd167)) &&(x > 10'd189) &&(x <10'd196) ) ||
    ( (y== ( 10'd168)) &&(x > 10'd189) &&(x <10'd195) ) ||
    ( (y== ( 10'd169)) &&(x > 10'd189) &&(x <10'd196) ) ||
    
    ( (x== ( 10'd290)) &&(y > 10'd37) &&(y <10'd50) )||//cloud3
    ( (x== ( 10'd291)) &&(y > 10'd37) &&(y <10'd50) ) ||
    ( (x== ( 10'd292)) &&(y > 10'd30) &&(y <10'd50) )||
    ( (x== ( 10'd293)) &&(y > 10'd37) &&(y <10'd50) ) ||
    ( (x== ( 10'd294)) &&(y > 10'd36) &&(y <10'd50) )||
    ( (x== ( 10'd295)) &&(y > 10'd37) &&(y <10'd50) ) ||
    ( (x== ( 10'd296)) &&(y > 10'd34) &&(y <10'd50) )||
    ( (x== ( 10'd297)) &&(y > 10'd33) &&(y <10'd50) ) ||
    ( (x== ( 10'd298)) &&(y > 10'd34) &&(y <10'd50) )||
    ( (x== ( 10'd299)) &&(y > 10'd32) &&(y <10'd50) ) ||
    ( (x== ( 10'd300)) &&(y > 10'd31) &&(y <10'd50) )||
    ( (x== ( 10'd301)) &&(y > 10'd32) &&(y <10'd50) ) ||
    ( (x== ( 10'd302)) &&(y > 10'd29) &&(y <10'd50) )||
    ( (x== ( 10'd303)) &&(y > 10'd28) &&(y <10'd50) ) ||
    ( (x== ( 10'd304)) &&(y > 10'd29) &&(y <10'd50) )||
    ( (x== ( 10'd305)) &&(y > 10'd28) &&(y <10'd50) ) ||
    ( (x== ( 10'd306)) &&(y > 10'd27) &&(y <10'd50) )||
    ( (x== ( 10'd307)) &&(y > 10'd28) &&(y <10'd50) ) ||
    ( (x== ( 10'd308)) &&(y > 10'd31) &&(y <10'd50) )||
    ( (x== ( 10'd309)) &&(y > 10'd30) &&(y <10'd50) ) ||
    ( (x== ( 10'd310)) &&(y > 10'd31) &&(y <10'd50) )||
    ( (x== ( 10'd311)) &&(y > 10'd32) &&(y <10'd50) ) ||
    ( (x== ( 10'd312)) &&(y > 10'd31) &&(y <10'd50) )||
    ( (x== ( 10'd313)) &&(y > 10'd32) &&(y <10'd50) ) ||
    ( (x== ( 10'd314)) &&(y > 10'd32) &&(y <10'd50) )||
    ( (x== ( 10'd315)) &&(y > 10'd35) &&(y <10'd50) ) ||
    ( (x== ( 10'd316)) &&(y > 10'd34) &&(y <10'd50) )||
    ( (x== ( 10'd317)) &&(y > 10'd35) &&(y <10'd50) ) ||
    ( (x== ( 10'd318)) &&(y > 10'd33) &&(y <10'd50) )||
    ( (x== ( 10'd319)) &&(y > 10'd33) &&(y <10'd50) ) ||
    ( (x== ( 10'd320)) &&(y > 10'd32) &&(y <10'd50) )||
    ( (x== ( 10'd321)) &&(y > 10'd33) &&(y <10'd50) ) ||
    ( (x== ( 10'd322)) &&(y > 10'd35) &&(y <10'd50) )||
    ( (x== ( 10'd323)) &&(y > 10'd34) &&(y <10'd50) ) ||
    ( (x== ( 10'd324)) &&(y > 10'd35) &&(y <10'd50) )||
    ( (x== ( 10'd325)) &&(y > 10'd36) &&(y <10'd50) ) ||
    ( (x== ( 10'd326)) &&(y > 10'd35) &&(y <10'd50) )||
    ( (x== ( 10'd327)) &&(y > 10'd36) &&(y <10'd50) ) ||
    ( (x== ( 10'd328)) &&(y > 10'd38) &&(y <10'd50) )||
    ( (x== ( 10'd329)) &&(y > 10'd37) &&(y <10'd50) ) ||
    ( (x== ( 10'd330)) &&(y > 10'd38) &&(y <10'd50) )||
    ( (x== ( 10'd331)) &&(y > 10'd37) &&(y <10'd50) ) ||
    ( (x== ( 10'd332)) &&(y > 10'd36) &&(y <10'd50) )||
    ( (x== ( 10'd333)) &&(y > 10'd37) &&(y <10'd50) ) ||
    ( (x== ( 10'd334)) &&(y > 10'd38) &&(y <10'd50) )||
    ( (x== ( 10'd335)) &&(y > 10'd37) &&(y <10'd50) ) ||
    ( (x== ( 10'd336)) &&(y > 10'd38) &&(y <10'd50) )||
    ( (x== ( 10'd337)) &&(y > 10'd36) &&(y <10'd50) ) ||
    ( (x== ( 10'd338)) &&(y > 10'd35) &&(y <10'd50) )||
    ( (x== ( 10'd339)) &&(y > 10'd35) &&(y <10'd50) ) ||
    ( (x== ( 10'd340)) &&(y > 10'd36) &&(y <10'd50) )||
    ( (x== ( 10'd341)) &&(y > 10'd33) &&(y <10'd50) ) ||
    ( (x== ( 10'd342)) &&(y > 10'd32) &&(y <10'd50) )||
    ( (x== ( 10'd343)) &&(y > 10'd33) &&(y <10'd50) ) ||
    ( (x== ( 10'd344)) &&(y > 10'd31) &&(y <10'd50) )||
    ( (x== ( 10'd345)) &&(y > 10'd30) &&(y <10'd50) ) ||
    ( (x== ( 10'd346)) &&(y > 10'd31) &&(y <10'd50) )||
    ( (x== ( 10'd347)) &&(y > 10'd29) &&(y <10'd50) ) ||
    ( (x== ( 10'd348)) &&(y > 10'd28) &&(y <10'd50) )||
    ( (x== ( 10'd349)) &&(y > 10'd29) &&(y <10'd50) ) ||
    ( (x== ( 10'd350)) &&(y > 10'd29) &&(y <10'd50) ) ||
    ( (y== ( 10'd41)) &&(x > 10'd286) &&(x <10'd290) ) ||//cloud3_left
    ( (y== ( 10'd42)) &&(x > 10'd285) &&(x <10'd290) ) ||
    ( (y== ( 10'd43)) &&(x > 10'd286) &&(x <10'd290) ) ||
    ( (y== ( 10'd44)) &&(x > 10'd285) &&(x <10'd290) ) ||
    ( (y== ( 10'd45)) &&(x > 10'd286) &&(x <10'd290) ) ||
    ( (y== ( 10'd46)) &&(x > 10'd285) &&(x <10'd290) ) ||
    ( (y== ( 10'd47)) &&(x > 10'd283) &&(x <10'd290) ) ||
    ( (y== ( 10'd48)) &&(x > 10'd284) &&(x <10'd290) ) ||
    ( (y== ( 10'd49)) &&(x > 10'd283) &&(x <10'd290) ) ||
    ( (y== ( 10'd30)) &&(x > 10'd350) &&(x <10'd352) ) ||//cloud3_right
    ( (y== ( 10'd31)) &&(x > 10'd350) &&(x <10'd351) ) ||
    ( (y== ( 10'd32)) &&(x > 10'd350) &&(x <10'd352) ) ||
    ( (y== ( 10'd33)) &&(x > 10'd350) &&(x <10'd353) ) ||
    ( (y== ( 10'd34)) &&(x > 10'd350) &&(x <10'd352) ) ||
    ( (y== ( 10'd35)) &&(x > 10'd350) &&(x <10'd353) ) ||
    ( (y== ( 10'd36)) &&(x > 10'd350) &&(x <10'd353) ) ||
    ( (y== ( 10'd37)) &&(x > 10'd350) &&(x <10'd354) ) ||
    ( (y== ( 10'd38)) &&(x > 10'd350) &&(x <10'd353) ) ||
    ( (y== ( 10'd39)) &&(x > 10'd350) &&(x <10'd354) ) ||
    ( (y== ( 10'd40)) &&(x > 10'd350) &&(x <10'd353) ) ||
    ( (y== ( 10'd41)) &&(x > 10'd350) &&(x <10'd353) ) ||
    ( (y== ( 10'd42)) &&(x > 10'd350) &&(x <10'd352) ) ||
    ( (y== ( 10'd43)) &&(x > 10'd350) &&(x <10'd353) ) ||
    ( (y== ( 10'd44)) &&(x > 10'd350) &&(x <10'd355) ) ||
    ( (y== ( 10'd45)) &&(x > 10'd350) &&(x <10'd354) ) ||
    ( (y== ( 10'd46)) &&(x > 10'd350) &&(x <10'd355) ) ||
    ( (y== ( 10'd47)) &&(x > 10'd350) &&(x <10'd356) ) ||
    ( (y== ( 10'd48)) &&(x > 10'd350) &&(x <10'd355) ) ||
    ( (y== ( 10'd49)) &&(x > 10'd350) &&(x <10'd356) ) ||
    ( (x== ( 10'd330)) &&(y > 10'd120) &&(y <10'd130) )||//cloud4
    ( (x== ( 10'd331)) &&(y > 10'd117) &&(y <10'd130) ) ||
    ( (x== ( 10'd332)) &&(y > 10'd116) &&(y <10'd130) )||
    ( (x== ( 10'd333)) &&(y > 10'd117) &&(y <10'd130) ) ||
    ( (x== ( 10'd334)) &&(y > 10'd116) &&(y <10'd130) )||
    ( (x== ( 10'd335)) &&(y > 10'd117) &&(y <10'd130) ) ||
    ( (x== ( 10'd336)) &&(y > 10'd114) &&(y <10'd130) )||
    ( (x== ( 10'd337)) &&(y > 10'd113) &&(y <10'd130) ) ||
    ( (x== ( 10'd338)) &&(y > 10'd114) &&(y <10'd130) )||
    ( (x== ( 10'd339)) &&(y > 10'd112) &&(y <10'd130) ) ||
    ( (x== ( 10'd340)) &&(y > 10'd111) &&(y <10'd130) )||
    ( (x== ( 10'd341)) &&(y > 10'd112) &&(y <10'd130) ) ||
    ( (x== ( 10'd342)) &&(y > 10'd113) &&(y <10'd130) )||
    ( (x== ( 10'd343)) &&(y > 10'd108) &&(y <10'd130) ) ||
    ( (x== ( 10'd344)) &&(y > 10'd109) &&(y <10'd130) )||
    ( (x== ( 10'd345)) &&(y > 10'd108) &&(y <10'd130) ) ||
    ( (x== ( 10'd346)) &&(y > 10'd107) &&(y <10'd130) )||
    ( (x== ( 10'd347)) &&(y > 10'd108) &&(y <10'd130) ) ||
    ( (x== ( 10'd348)) &&(y > 10'd111) &&(y <10'd130) )||
    ( (x== ( 10'd349)) &&(y > 10'd110) &&(y <10'd130) ) ||
    ( (x== ( 10'd350)) &&(y > 10'd111) &&(y <10'd130) )||
    ( (x== ( 10'd351)) &&(y > 10'd112) &&(y <10'd130) ) ||
    ( (x== ( 10'd352)) &&(y > 10'd111) &&(y <10'd130) )||
    ( (x== ( 10'd353)) &&(y > 10'd112) &&(y <10'd130) ) ||
    ( (x== ( 10'd354)) &&(y > 10'd112) &&(y <10'd130) )||
    ( (x== ( 10'd355)) &&(y > 10'd115) &&(y <10'd130) ) ||
    ( (x== ( 10'd356)) &&(y > 10'd114) &&(y <10'd130) )||
    ( (x== ( 10'd357)) &&(y > 10'd115) &&(y <10'd130) ) ||
    ( (x== ( 10'd358)) &&(y > 10'd113) &&(y <10'd130) )||
    ( (x== ( 10'd359)) &&(y > 10'd113) &&(y <10'd130) ) ||
    ( (x== ( 10'd360)) &&(y > 10'd112) &&(y <10'd130) )||
    ( (x== ( 10'd361)) &&(y > 10'd113) &&(y <10'd130) ) ||
    ( (x== ( 10'd362)) &&(y > 10'd115) &&(y <10'd130) )||
    ( (x== ( 10'd363)) &&(y > 10'd114) &&(y <10'd130) ) ||
    ( (x== ( 10'd364)) &&(y > 10'd115) &&(y <10'd130) )||
    ( (x== ( 10'd365)) &&(y > 10'd116) &&(y <10'd130) ) ||
    ( (x== ( 10'd366)) &&(y > 10'd115) &&(y <10'd130) )||
    ( (x== ( 10'd367)) &&(y > 10'd116) &&(y <10'd130) ) ||
    ( (x== ( 10'd368)) &&(y > 10'd118) &&(y <10'd130) )||
    ( (x== ( 10'd369)) &&(y > 10'd117) &&(y <10'd130) ) ||
    
    ( (y== ( 10'd121)) &&(x > 10'd326) &&(x <10'd330) ) ||//cloud4_left
    ( (y== ( 10'd122)) &&(x > 10'd325) &&(x <10'd330) ) ||
    ( (y== ( 10'd123)) &&(x > 10'd326) &&(x <10'd330) ) ||
    ( (y== ( 10'd124)) &&(x > 10'd325) &&(x <10'd330) ) ||
    ( (y== ( 10'd125)) &&(x > 10'd326) &&(x <10'd330) ) ||
    ( (y== ( 10'd126)) &&(x > 10'd325) &&(x <10'd330) ) ||
    ( (y== ( 10'd127)) &&(x > 10'd323) &&(x <10'd330) ) ||
    ( (y== ( 10'd128)) &&(x > 10'd324) &&(x <10'd330) ) ||
    ( (y== ( 10'd129)) &&(x > 10'd323) &&(x <10'd330) ) ||
    ( (y== ( 10'd118)) &&(x > 10'd369) &&(x <10'd371) ) ||//cloud4_right
    ( (y== ( 10'd119)) &&(x > 10'd369) &&(x <10'd370) ) ||
    ( (y== ( 10'd120)) &&(x > 10'd369) &&(x <10'd371) ) ||
    ( (y== ( 10'd121)) &&(x > 10'd369) &&(x <10'd372) ) ||
    ( (y== ( 10'd122)) &&(x > 10'd369) &&(x <10'd371) ) ||
    ( (y== ( 10'd123)) &&(x > 10'd369) &&(x <10'd372) ) ||
    ( (y== ( 10'd124)) &&(x > 10'd369) &&(x <10'd372) ) ||
    ( (y== ( 10'd125)) &&(x > 10'd369) &&(x <10'd373) ) ||
    ( (y== ( 10'd126)) &&(x > 10'd369) &&(x <10'd372) ) ||
    ( (y== ( 10'd127)) &&(x > 10'd369) &&(x <10'd373) ) ||
    ( (y== ( 10'd128)) &&(x > 10'd369) &&(x <10'd372) ) ||
    ( (y== ( 10'd129)) &&(x > 10'd369) &&(x <10'd372) ) ||
    ( (x== ( 10'd440)) &&(y > 10'd97) &&(y <10'd110) )||//cloud5
    ( (x== ( 10'd441)) &&(y > 10'd97) &&(y <10'd110) ) ||
    ( (x== ( 10'd442)) &&(y > 10'd90) &&(y <10'd110) )||
    ( (x== ( 10'd443)) &&(y > 10'd97) &&(y <10'd110) ) ||
    ( (x== ( 10'd444)) &&(y > 10'd96) &&(y <10'd110) )||
    ( (x== ( 10'd445)) &&(y > 10'd97) &&(y <10'd110) ) ||
    ( (x== ( 10'd446)) &&(y > 10'd94) &&(y <10'd110) )||
    ( (x== ( 10'd447)) &&(y > 10'd93) &&(y <10'd110) ) ||
    ( (x== ( 10'd448)) &&(y > 10'd94) &&(y <10'd110) )||
    ( (x== ( 10'd449)) &&(y > 10'd92) &&(y <10'd110) ) ||
    ( (x== ( 10'd450)) &&(y > 10'd91) &&(y <10'd110) )||
    ( (x== ( 10'd451)) &&(y > 10'd92) &&(y <10'd110) ) ||
    ( (x== ( 10'd452)) &&(y > 10'd89) &&(y <10'd110) )||
    ( (x== ( 10'd453)) &&(y > 10'd88) &&(y <10'd110) ) ||
    ( (x== ( 10'd454)) &&(y > 10'd89) &&(y <10'd110) )||
    ( (x== ( 10'd455)) &&(y > 10'd88) &&(y <10'd110) ) ||
    ( (x== ( 10'd456)) &&(y > 10'd87) &&(y <10'd110) )||
    ( (x== ( 10'd457)) &&(y > 10'd88) &&(y <10'd110) ) ||
    ( (x== ( 10'd458)) &&(y > 10'd91) &&(y <10'd110) )||
    ( (x== ( 10'd459)) &&(y > 10'd90) &&(y <10'd110) ) ||
    ( (x== ( 10'd460)) &&(y > 10'd91) &&(y <10'd110) )||
    ( (x== ( 10'd461)) &&(y > 10'd92) &&(y <10'd110) ) ||
    ( (x== ( 10'd462)) &&(y > 10'd91) &&(y <10'd110) )||
    ( (x== ( 10'd463)) &&(y > 10'd92) &&(y <10'd110) ) ||
    ( (x== ( 10'd464)) &&(y > 10'd92) &&(y <10'd110) )||
    ( (x== ( 10'd465)) &&(y > 10'd95) &&(y <10'd110) ) ||
    ( (x== ( 10'd466)) &&(y > 10'd94) &&(y <10'd110) )||
    ( (x== ( 10'd467)) &&(y > 10'd95) &&(y <10'd110) ) ||
    ( (x== ( 10'd468)) &&(y > 10'd93) &&(y <10'd110) )||
    ( (x== ( 10'd469)) &&(y > 10'd93) &&(y <10'd110) ) ||
    ( (x== ( 10'd470)) &&(y > 10'd92) &&(y <10'd110) )||
    ( (x== ( 10'd471)) &&(y > 10'd93) &&(y <10'd110) ) ||
    ( (x== ( 10'd472)) &&(y > 10'd95) &&(y <10'd110) )||
    ( (x== ( 10'd473)) &&(y > 10'd94) &&(y <10'd110) ) ||
    ( (x== ( 10'd474)) &&(y > 10'd95) &&(y <10'd110) )||
    ( (x== ( 10'd475)) &&(y > 10'd96) &&(y <10'd110) ) ||
    ( (x== ( 10'd476)) &&(y > 10'd95) &&(y <10'd110) )||
    ( (x== ( 10'd477)) &&(y > 10'd96) &&(y <10'd110) ) ||
    ( (x== ( 10'd478)) &&(y > 10'd98) &&(y <10'd110) )||
    ( (x== ( 10'd479)) &&(y > 10'd97) &&(y <10'd110) ) ||
    ( (x== ( 10'd480)) &&(y > 10'd98) &&(y <10'd110) )||
    ( (x== ( 10'd481)) &&(y > 10'd97) &&(y <10'd110) ) ||
    ( (x== ( 10'd482)) &&(y > 10'd96) &&(y <10'd110) )||
    ( (x== ( 10'd483)) &&(y > 10'd97) &&(y <10'd110) ) ||
    ( (x== ( 10'd484)) &&(y > 10'd98) &&(y <10'd110) )||
    ( (x== ( 10'd485)) &&(y > 10'd97) &&(y <10'd110) ) ||
    ( (x== ( 10'd486)) &&(y > 10'd98) &&(y <10'd110) )||
    ( (x== ( 10'd487)) &&(y > 10'd96) &&(y <10'd110) ) ||
    ( (x== ( 10'd488)) &&(y > 10'd95) &&(y <10'd110) )||
    ( (x== ( 10'd489)) &&(y > 10'd95) &&(y <10'd110) ) ||
    ( (x== ( 10'd490)) &&(y > 10'd96) &&(y <10'd110) )||
    ( (x== ( 10'd491)) &&(y > 10'd93) &&(y <10'd110) ) ||
    ( (x== ( 10'd492)) &&(y > 10'd92) &&(y <10'd110) )||
    ( (x== ( 10'd493)) &&(y > 10'd93) &&(y <10'd110) ) ||
    ( (x== ( 10'd494)) &&(y > 10'd91) &&(y <10'd110) )||
    ( (x== ( 10'd495)) &&(y > 10'd90) &&(y <10'd110) ) ||
    ( (x== ( 10'd496)) &&(y > 10'd91) &&(y <10'd110) )||
    ( (x== ( 10'd497)) &&(y > 10'd89) &&(y <10'd110) ) ||
    ( (x== ( 10'd498)) &&(y > 10'd88) &&(y <10'd110) )||
    ( (x== ( 10'd499)) &&(y > 10'd89) &&(y <10'd110) ) ||
    ( (x== ( 10'd500)) &&(y > 10'd89) &&(y <10'd110) ) ||
    ( (y== ( 10'd101)) &&(x > 10'd436) &&(x <10'd440) ) ||//cloud5_left
    ( (y== ( 10'd102)) &&(x > 10'd435) &&(x <10'd440) ) ||
    ( (y== ( 10'd103)) &&(x > 10'd436) &&(x <10'd440) ) ||
    ( (y== ( 10'd104)) &&(x > 10'd435) &&(x <10'd440) ) ||
    ( (y== ( 10'd105)) &&(x > 10'd436) &&(x <10'd440) ) ||
    ( (y== ( 10'd106)) &&(x > 10'd435) &&(x <10'd440) ) ||
    ( (y== ( 10'd107)) &&(x > 10'd433) &&(x <10'd440) ) ||
    ( (y== ( 10'd108)) &&(x > 10'd434) &&(x <10'd440) ) ||
    ( (y== ( 10'd109)) &&(x > 10'd433) &&(x <10'd440) ) ||
    ( (y== ( 10'd90)) &&(x > 10'd500) &&(x <10'd502) ) ||//cloud5_right
    ( (y== ( 10'd91)) &&(x > 10'd500) &&(x <10'd501) ) ||
    ( (y== ( 10'd92)) &&(x > 10'd500) &&(x <10'd502) ) ||
    ( (y== ( 10'd93)) &&(x > 10'd500) &&(x <10'd503) ) ||
    ( (y== ( 10'd94)) &&(x > 10'd500) &&(x <10'd502) ) ||
    ( (y== ( 10'd95)) &&(x > 10'd500) &&(x <10'd503) ) ||
    ( (y== ( 10'd96)) &&(x > 10'd500) &&(x <10'd503) ) ||
    ( (y== ( 10'd97)) &&(x > 10'd500) &&(x <10'd504) ) ||
    ( (y== ( 10'd98)) &&(x > 10'd500) &&(x <10'd503) ) ||
    ( (y== ( 10'd99)) &&(x > 10'd500) &&(x <10'd504) ) ||
    ( (y== ( 10'd100)) &&(x > 10'd500) &&(x <10'd503) ) ||
    ( (y== ( 10'd101)) &&(x > 10'd500) &&(x <10'd503) ) ||
    ( (y== ( 10'd102)) &&(x > 10'd500) &&(x <10'd502) ) ||
    ( (y== ( 10'd103)) &&(x > 10'd500) &&(x <10'd503) ) ||
    ( (y== ( 10'd104)) &&(x > 10'd500) &&(x <10'd505) ) ||
    ( (y== ( 10'd105)) &&(x > 10'd500) &&(x <10'd504) ) ||
    ( (y== ( 10'd106)) &&(x > 10'd500) &&(x <10'd505) ) ||
    ( (y== ( 10'd107)) &&(x > 10'd500) &&(x <10'd506) ) ||
    ( (y== ( 10'd108)) &&(x > 10'd500) &&(x <10'd505) ) ||
    ( (y== ( 10'd109)) &&(x > 10'd500) &&(x <10'd506) ) 
    
    
    
    ;
    assign sun =
    ( (x>= ( 10'd565)) &&(x<= ( 10'd605)) &&(y >= 10'd55) &&(y <=10'd95) ) ||
    ( (x>= ( 10'd583)) &&(x<= ( 10'd587)) &&(y >= 10'd98) &&(y <=10'd110) ) ||//6
    ( (x>= ( 10'd583)) &&(x<= ( 10'd587)) &&(y >= 10'd40) &&(y <=10'd52) ) ||//2
    ( (x>= ( 10'd550)) &&(x<= ( 10'd562)) &&(y >= 10'd73) &&(y <=10'd77) ) ||//8
    ( (x>= ( 10'd608)) &&(x<= ( 10'd620)) &&(y >= 10'd73) &&(y <=10'd77) )  ||//4
    ( (x== ( 10'd562)) &&(y > 10'd96) &&(y <10'd104) )||//7
    ( (x== ( 10'd561)) &&(y > 10'd97) &&(y <10'd105) )||
    ( (x== ( 10'd560)) &&(y > 10'd98) &&(y <10'd106) )||
    ( (x== ( 10'd559)) &&(y > 10'd99) &&(y <10'd107) )||
    ( (x== ( 10'd558)) &&(y > 10'd100) &&(y <10'd108) )||
    ( (x== ( 10'd557)) &&(y > 10'd101) &&(y <10'd109) )||
    ( (x== ( 10'd556)) &&(y > 10'd102) &&(y <10'd110) ) ||
    ( (x== ( 10'd555)) &&(y > 10'd103) &&(y <10'd111) ) ||
    ( (x== ( 10'd554)) &&(y > 10'd104) &&(y <10'd112) ) ||
    ( (x== ( 10'd562)) &&(y > 10'd44) &&(y <10'd52) )||//1
    ( (x== ( 10'd561)) &&(y > 10'd43) &&(y <10'd51) )||
    ( (x== ( 10'd560)) &&(y > 10'd42) &&(y <10'd50) )||
    ( (x== ( 10'd559)) &&(y > 10'd41) &&(y <10'd49) )||
    ( (x== ( 10'd558)) &&(y > 10'd40) &&(y <10'd48) )||
    ( (x== ( 10'd557)) &&(y > 10'd39) &&(y <10'd47) )||
    ( (x== ( 10'd556)) &&(y > 10'd38) &&(y <10'd46) ) ||
    ( (x== ( 10'd555)) &&(y > 10'd37) &&(y <10'd45) ) ||
    ( (x== ( 10'd554)) &&(y > 10'd36) &&(y <10'd44) ) ||
    ( (x== ( 10'd608)) &&(y > 10'd44) &&(y <10'd52) )||//3
    ( (x== ( 10'd609)) &&(y > 10'd43) &&(y <10'd51) )||
    ( (x== ( 10'd610)) &&(y > 10'd42) &&(y <10'd50) )||
    ( (x== ( 10'd611)) &&(y > 10'd41) &&(y <10'd49) )||
    ( (x== ( 10'd612)) &&(y > 10'd40) &&(y <10'd48) )||
    ( (x== ( 10'd613)) &&(y > 10'd39) &&(y <10'd47) )||
    ( (x== ( 10'd614)) &&(y > 10'd38) &&(y <10'd46) ) ||
    ( (x== ( 10'd615)) &&(y > 10'd37) &&(y <10'd45) ) ||
    ( (x== ( 10'd616)) &&(y > 10'd36) &&(y <10'd44) ) ||
    ( (x== ( 10'd608)) &&(y > 10'd96) &&(y <10'd104) )||//5
    ( (x== ( 10'd609)) &&(y > 10'd97) &&(y <10'd105) )||
    ( (x== ( 10'd610)) &&(y > 10'd98) &&(y <10'd106) )||
    ( (x== ( 10'd611)) &&(y > 10'd99) &&(y <10'd107) )||
    ( (x== ( 10'd612)) &&(y > 10'd100) &&(y <10'd108) )||
    ( (x== ( 10'd613)) &&(y > 10'd101) &&(y <10'd109) )||
    ( (x== ( 10'd614)) &&(y > 10'd102) &&(y <10'd110) ) ||
    ( (x== ( 10'd615)) &&(y > 10'd103) &&(y <10'd111) ) ||
    ( (x== ( 10'd616)) &&(y > 10'd104) &&(y <10'd112) ) 
    ;   
    assign dino_draw =  
    ( (x== (dino_x + 10'd3)) &&(y > (dino_y+10'd35)) &&(y <dino_y+10'd55) )||
    ( (x== (dino_x + 10'd4)) &&(y > (dino_y+10'd38)) &&(y <dino_y+10'd58) )||
    ( (x== (dino_x + 10'd5)) &&(y > (dino_y+10'd41)) &&(y <dino_y+10'd61) )||
    ( (x== (dino_x + 10'd6)) &&(y > (dino_y+10'd44)) &&(y <dino_y+10'd61) )||
    ( (x== (dino_x + 10'd7)) &&(y > (dino_y+10'd44)) &&(y <dino_y+10'd61) )||
    ( (x== (dino_x + 10'd8)) &&(y > (dino_y+10'd44)) &&(y <dino_y+10'd71) )||
    ( (x== (dino_x + 10'd9)) &&(y > (dino_y+10'd41)) &&(y <dino_y+10'd79) )||
    ( (x== (dino_x + 10'd10)) &&(y > (dino_y+10'd38)) &&(y <dino_y+10'd75) )||
    ( (x== (dino_x + 10'd10)) &&(y > (dino_y+10'd77)) &&(y <dino_y+10'd79) )||
    ( (x== (dino_x + 10'd11)) &&(y > (dino_y+10'd35)) &&(y <dino_y+10'd72) )||
    ( (x== (dino_x + 10'd12)) &&(y > (dino_y+10'd35)) &&(y <dino_y+10'd72) )||
    ( (x== (dino_x + 10'd13)) &&(y > (dino_y+10'd32)) &&(y <dino_y+10'd69) )||
    ( (x== (dino_x + 10'd14)) &&(y > (dino_y+10'd32)) &&(y <dino_y+10'd69) )||
    ( (x== (dino_x + 10'd15)) &&(y > (dino_y+10'd29)) &&(y <dino_y+10'd72) )||
    ( (x== (dino_x + 10'd16)) &&(y > (dino_y+10'd29)) &&(y <dino_y+10'd72) )||
    ( (x== (dino_x + 10'd17)) &&(y > (dino_y+10'd29)) &&(y <dino_y+10'd72) )||
    ( (x== (dino_x + 10'd17)) &&(y > (dino_y+10'd44)) &&(y <dino_y+10'd61) )||
    ( (x== (dino_x + 10'd18)) &&(y > (dino_y+10'd44)) &&(y <dino_y+10'd71) )||
    ( (x== (dino_x + 10'd18)) &&(y > (dino_y+10'd29)) &&(y <dino_y+10'd72) )||
    ( (x== (dino_x + 10'd19)) &&(y > (dino_y+10'd41)) &&(y <dino_y+10'd79) )||
    ( (x== (dino_x + 10'd19)) &&(y > (dino_y+10'd29)) &&(y <dino_y+10'd72) )||
    ( (x== (dino_x + 10'd20)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd60) )||
    ( (x== (dino_x + 10'd20)) &&(y > (dino_y+10'd77)) &&(y <dino_y+10'd79) )||
    ( (x== (dino_x + 10'd21)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd3) )||
    ( (x== (dino_x + 10'd21)) &&(y > (dino_y+10'd5)) &&(y <dino_y+10'd57) )||
    ( (x== (dino_x + 10'd22)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd3) )||
    ( (x== (dino_x + 10'd22)) &&(y > (dino_y+10'd5)) &&(y <dino_y+10'd57) )||
    ( (x== (dino_x + 10'd23)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd54) )||
    ( (x== (dino_x + 10'd24)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd24)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd24)) &&(y > (dino_y+10'd34)) &&(y <dino_y+10'd37) )||
    ( (x== (dino_x + 10'd25)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd25)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd25)) &&(y > (dino_y+10'd34)) &&(y <dino_y+10'd37) )||
    ( (x== (dino_x + 10'd26)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd26)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd26)) &&(y > (dino_y+10'd34)) &&(y <dino_y+10'd40) )||
    ( (x== (dino_x + 10'd27)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd27)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd27)) &&(y > (dino_y+10'd35)) &&(y <dino_y+10'd40) )||
    ( (x== (dino_x + 10'd28)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd28)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd29)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd29)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd30)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd30)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd31)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd31)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd32)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd32)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd33)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd33)) &&(y > (dino_y+10'd27)) &&(y <dino_y+10'd30) )||
    ( (x== (dino_x + 10'd34)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd35)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd36)) &&(y > (dino_y+10'd1)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd37)) &&(y > (dino_y+10'd4)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd38)) &&(y > (dino_y+10'd4)) &&(y <dino_y+10'd27) )||
    ( (x== (dino_x + 10'd39)) &&(y > (dino_y+10'd4)) &&(y <dino_y+10'd27) )
    ;
    assign obtacle_draw =  
    ( (x== (obtacle_x + 10'd2)) &&(y > (obtacle_y+10'd15)) &&(y <obtacle_y+10'd36) )||
    ( (x== (obtacle_x + 10'd3)) &&(y > (obtacle_y+10'd14)) &&(y <obtacle_y+10'd36) )||
    ( (x== (obtacle_x + 10'd4)) &&(y > (obtacle_y+10'd15)) &&(y <obtacle_y+10'd36) )||
    ( (x== (obtacle_x + 10'd5)) &&(y > (obtacle_y+10'd33)) &&(y <obtacle_y+10'd36) )||
    ( (x== (obtacle_x + 10'd6)) &&(y > (obtacle_y+10'd33)) &&(y <obtacle_y+10'd36) )||
    ( (x== (obtacle_x + 10'd7)) &&(y > (obtacle_y+10'd3)) &&(y <obtacle_y+10'd50) )||
    ( (x== (obtacle_x + 10'd8)) &&(y > (obtacle_y+10'd2)) &&(y <obtacle_y+10'd50) )||
    ( (x== (obtacle_x + 10'd9)) &&(y > (obtacle_y+10'd2)) &&(y <obtacle_y+10'd50) )||
    ( (x== (obtacle_x + 10'd10)) &&(y > (obtacle_y+10'd3)) &&(y <obtacle_y+10'd50) )||
    ( (x== (obtacle_x + 10'd11)) &&(y > (obtacle_y+10'd32)) &&(y <obtacle_y+10'd35) )||
    ( (x== (obtacle_x + 10'd12)) &&(y > (obtacle_y+10'd32)) &&(y <obtacle_y+10'd35) )||
    ( (x== (obtacle_x + 10'd13)) &&(y > (obtacle_y+10'd10)) &&(y <obtacle_y+10'd35) )||
    ( (x== (obtacle_x + 10'd14)) &&(y > (obtacle_y+10'd9)) &&(y <obtacle_y+10'd35) )||
    ( (x== (obtacle_x + 10'd15)) &&(y > (obtacle_y+10'd10)) &&(y <obtacle_y+10'd35) )||
    ( (x== (obtacle_x + 10'd17)) &&(y > (obtacle_y+10'd9)) &&(y <obtacle_y+10'd38) )||
    ( (x== (obtacle_x + 10'd18)) &&(y > (obtacle_y+10'd8)) &&(y <obtacle_y+10'd38) )||
    ( (x== (obtacle_x + 10'd19)) &&(y > (obtacle_y+10'd9)) &&(y <obtacle_y+10'd38) )||
    ( (x== (obtacle_x + 10'd20)) &&(y > (obtacle_y+10'd35)) &&(y <obtacle_y+10'd38) )||
    ( (x== (obtacle_x + 10'd21)) &&(y > (obtacle_y+10'd35)) &&(y <obtacle_y+10'd38) )||
    ( (x== (obtacle_x + 10'd22)) &&(y > (obtacle_y+10'd3)) &&(y <obtacle_y+10'd50) )||
    ( (x== (obtacle_x + 10'd23)) &&(y > (obtacle_y+10'd2)) &&(y <obtacle_y+10'd50) )||
    ( (x== (obtacle_x + 10'd24)) &&(y > (obtacle_y+10'd2)) &&(y <obtacle_y+10'd50) )||
    ( (x== (obtacle_x + 10'd25)) &&(y > (obtacle_y+10'd3)) &&(y <obtacle_y+10'd50) )||
    ( (x== (obtacle_x + 10'd26)) &&(y > (obtacle_y+10'd32)) &&(y <obtacle_y+10'd35) )||
    ( (x== (obtacle_x + 10'd27)) &&(y > (obtacle_y+10'd32)) &&(y <obtacle_y+10'd35) )||
    ( (x== (obtacle_x + 10'd28)) &&(y > (obtacle_y+10'd32)) &&(y <obtacle_y+10'd45) )||
    ( (x== (obtacle_x + 10'd29)) &&(y > (obtacle_y+10'd32)) &&(y <obtacle_y+10'd45) )
    ;
    assign black =
    ( (x== 10'd70) &&(y > 10'd415) &&(y <10'd435) )|| //dino1
    ( (x== 10'd71) &&(y > 10'd418) &&(y <10'd438) )||
    ( (x== 10'd72) &&(y > 10'd421) &&(y <10'd441 ))||
    ( (x== 10'd73) &&(y > 10'd424) &&(y <10'd441 ))||
    ( (x== 10'd74) &&(y > 10'd424) &&(y <10'd441 ))||
    ( (x== 10'd75) &&(y > 10'd424) &&(y <10'd451 ))||
    ( (x== 10'd76) &&(y > 10'd421) &&(y <10'd459 ))||
    ( (x== 10'd77) &&(y > 10'd418) &&(y <10'd455 ))||
    ( (x== 10'd77) &&(y > 10'd457) &&(y <10'd459 ))||
    ( (x== 10'd78) &&(y > 10'd415) &&(y <10'd452) )||
    ( (x== 10'd79) &&(y > 10'd415) &&(y <10'd452) )||
    ( (x== 10'd80) &&(y > 10'd412) &&(y <10'd449) )||
    ( (x==  10'd81) &&(y > 10'd412) &&(y <10'd449) )||
    ( (x==  10'd82) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x==  10'd83) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x== 10'd84) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x== 10'd84) &&(y > 10'd424) &&(y <10'd441) )||
    ( (x==  10'd85) &&(y > 10'd424) &&(y <10'd451) )||
    ( (x==  10'd85) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x==  10'd86) &&(y > 10'd421) &&(y <10'd459) )||
    ( (x==  10'd86) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x==  10'd87) &&(y > 10'd381) &&(y <10'd440) )||
    ( (x== 10'd87) &&(y > 10'd457) &&(y <10'd459) )||
    ( (x==  10'd88) &&(y > 10'd381) &&(y <10'd383) )||
    ( (x==  10'd88) &&(y > 10'd385) &&(y <10'd437) )||
    ( (x==  10'd89) &&(y > 10'd381) &&(y <10'd383) )||
    ( (x==  10'd89) &&(y > 10'd385) &&(y <10'd437) )||
    ( (x==  10'd90) &&(y > 10'd381) &&(y <10'd434) )||
    ( (x==  10'd91) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd91) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd91) &&(y > 10'd414) &&(y <10'd417) )||
    ( (x==  10'd92) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd92) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd92) &&(y > 10'd414) &&(y <10'd417) )||
    ( (x==  10'd93) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd93) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x== 10'd93) &&(y > 10'd414) &&(y <10'd420) )||
    ( (x==   10'd94) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd94) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x== 10'd94) &&(y > 10'd415) &&(y <10'd420) )||
    ( (x==  10'd95) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd95) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==   10'd96) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd96) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd97) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==   10'd97) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==   10'd98) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==   10'd98) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==   10'd99) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd99) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd100) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==   10'd100) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd101) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd102) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd103) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==   10'd104) &&(y > 10'd384) &&(y <10'd407) )||
    ( (x==   10'd105) &&(y > 10'd384) &&(y <10'd407) )||
    ( (x==   10'd106) &&(y > 10'd384) &&(y <10'd407) ) ||
    ( (x== 10'd198) &&(y > 10'd355) &&(y <10'd375) )|| //dino2
    ( (x== 10'd199) &&(y > 10'd358) &&(y <10'd378) )||
    ( (x== 10'd200) &&(y > 10'd361) &&(y <10'd381 ))||
    ( (x== 10'd201) &&(y > 10'd364) &&(y <10'd381 ))||
    ( (x== 10'd202) &&(y > 10'd364) &&(y <10'd381 ))||
    ( (x== 10'd203) &&(y > 10'd364) &&(y <10'd391 ))||
    ( (x== 10'd204) &&(y > 10'd361) &&(y <10'd399 ))||
    ( (x== 10'd205) &&(y > 10'd358) &&(y <10'd395 ))||
    ( (x== 10'd205) &&(y > 10'd397) &&(y <10'd399 ))||
    ( (x== 10'd206) &&(y > 10'd355) &&(y <10'd392) )||
    ( (x== 10'd207) &&(y > 10'd355) &&(y <10'd392) )||
    ( (x== 10'd208) &&(y > 10'd352) &&(y <10'd389) )||
    ( (x==  10'd209) &&(y > 10'd352) &&(y <10'd389) )||
    ( (x==  10'd210) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x==  10'd211) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x== 10'd212) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x== 10'd212) &&(y > 10'd364) &&(y <10'd381) )||
    ( (x==  10'd213) &&(y > 10'd364) &&(y <10'd391) )||
    ( (x==  10'd213) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x==  10'd214) &&(y > 10'd361) &&(y <10'd399) )||
    ( (x==  10'd214) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x==  10'd215) &&(y > 10'd321) &&(y <10'd380) )||
    ( (x== 10'd215) &&(y > 10'd397) &&(y <10'd399) )||
    ( (x==  10'd216) &&(y > 10'd321) &&(y <10'd323) )||
    ( (x==  10'd216) &&(y > 10'd325) &&(y <10'd377) )||
    ( (x==  10'd217) &&(y > 10'd321) &&(y <10'd323) )||
    ( (x==  10'd217) &&(y > 10'd325) &&(y <10'd377) )||
    ( (x==  10'd218) &&(y > 10'd321) &&(y <10'd374) )||
    ( (x==  10'd219) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd219) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd219) &&(y > 10'd354) &&(y <10'd357) )||
    ( (x==  10'd220) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd220) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd220) &&(y > 10'd354) &&(y <10'd357) )||
    ( (x==  10'd221) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd221) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x== 10'd221) &&(y > 10'd354) &&(y <10'd360) )||
    ( (x==   10'd222) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd222) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x== 10'd222) &&(y > 10'd355) &&(y <10'd360) )||
    ( (x==  10'd223) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd223) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==   10'd224) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd224) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd225) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==   10'd225) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==   10'd226) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==   10'd226) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==   10'd227) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd227) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd228) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==   10'd228) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd229) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd230) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd231) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==   10'd232) &&(y > 10'd324) &&(y <10'd347) )||
    ( (x==   10'd233) &&(y > 10'd324) &&(y <10'd347) )||
    ( (x==   10'd234) &&(y > 10'd324) &&(y <10'd347) ) ||
    ( (x== 10'd326) &&(y > 10'd295) &&(y <10'd315) )|| //dino3
    ( (x== 10'd327) &&(y > 10'd298) &&(y <10'd318) )||
    ( (x== 10'd328) &&(y > 10'd301) &&(y <10'd321 ))||
    ( (x== 10'd329) &&(y > 10'd304) &&(y <10'd321 ))||
    ( (x== 10'd330) &&(y > 10'd304) &&(y <10'd321 ))||
    ( (x== 10'd331) &&(y > 10'd304) &&(y <10'd331 ))||
    ( (x== 10'd332) &&(y > 10'd301) &&(y <10'd339 ))||
    ( (x== 10'd333) &&(y > 10'd298) &&(y <10'd335 ))||
    ( (x== 10'd333) &&(y > 10'd337) &&(y <10'd339 ))||
    ( (x== 10'd334) &&(y > 10'd295) &&(y <10'd332) )||
    ( (x== 10'd335) &&(y > 10'd295) &&(y <10'd332) )||
    ( (x== 10'd336) &&(y > 10'd292) &&(y <10'd329) )||
    ( (x==  10'd337) &&(y > 10'd292) &&(y <10'd329) )||
    ( (x==  10'd338) &&(y > 10'd289) &&(y <10'd332) )||
    ( (x==  10'd339) &&(y > 10'd289) &&(y <10'd332) )||
    ( (x== 10'd340) &&(y > 10'd289) &&(y <10'd332) )||
    ( (x== 10'd340) &&(y > 10'd304) &&(y <10'd321) )||
    ( (x==  10'd341) &&(y > 10'd304) &&(y <10'd331) )||
    ( (x==  10'd341) &&(y > 10'd289) &&(y <10'd332) )||
    ( (x==  10'd342) &&(y > 10'd301) &&(y <10'd339) )||
    ( (x==  10'd342) &&(y > 10'd289) &&(y <10'd332) )||
    ( (x==  10'd343) &&(y > 10'd261) &&(y <10'd320) )||
    ( (x== 10'd343) &&(y > 10'd337) &&(y <10'd339) )||
    ( (x==  10'd344) &&(y > 10'd261) &&(y <10'd263) )||
    ( (x==  10'd344) &&(y > 10'd265) &&(y <10'd317) )||
    ( (x==  10'd345) &&(y > 10'd261) &&(y <10'd263) )||
    ( (x==  10'd345) &&(y > 10'd265) &&(y <10'd317) )||
    ( (x==  10'd346) &&(y > 10'd261) &&(y <10'd314) )||
    ( (x==  10'd347) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd347) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x==  10'd347) &&(y > 10'd294) &&(y <10'd297) )||
    ( (x==  10'd348) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd348) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x==  10'd348) &&(y > 10'd294) &&(y <10'd297) )||
    ( (x==  10'd349) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd349) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x== 10'd349) &&(y > 10'd294) &&(y <10'd300) )||
    ( (x==   10'd350) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd350) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x== 10'd350) &&(y > 10'd295) &&(y <10'd300) )||
    ( (x==  10'd351) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd351) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x==   10'd352) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd352) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x==  10'd353) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==   10'd353) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x==   10'd354) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==   10'd354) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x==   10'd355) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd355) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x==  10'd356) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==   10'd356) &&(y > 10'd287) &&(y <10'd290) )||
    ( (x==  10'd357) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd358) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==  10'd359) &&(y > 10'd261) &&(y <10'd287) )||
    ( (x==   10'd360) &&(y > 10'd264) &&(y <10'd287) )||
    ( (x==   10'd361) &&(y > 10'd264) &&(y <10'd287) )||
    ( (x==   10'd362) &&(y > 10'd264) &&(y <10'd287) ) ||
    ( (x== 10'd454) &&(y > 10'd355) &&(y <10'd375) )|| //dino4
    ( (x== 10'd455) &&(y > 10'd358) &&(y <10'd378) )||
    ( (x== 10'd456) &&(y > 10'd361) &&(y <10'd381 ))||
    ( (x== 10'd457) &&(y > 10'd364) &&(y <10'd381 ))||
    ( (x== 10'd458) &&(y > 10'd364) &&(y <10'd381 ))||
    ( (x== 10'd459) &&(y > 10'd364) &&(y <10'd391 ))||
    ( (x== 10'd460) &&(y > 10'd361) &&(y <10'd399 ))||
    ( (x== 10'd461) &&(y > 10'd358) &&(y <10'd395 ))||
    ( (x== 10'd461) &&(y > 10'd397) &&(y <10'd399 ))||
    ( (x== 10'd462) &&(y > 10'd355) &&(y <10'd392) )||
    ( (x== 10'd463) &&(y > 10'd355) &&(y <10'd392) )||
    ( (x== 10'd464) &&(y > 10'd352) &&(y <10'd389) )||
    ( (x==  10'd465) &&(y > 10'd352) &&(y <10'd389) )||
    ( (x==  10'd466) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x==  10'd467) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x== 10'd468) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x== 10'd468) &&(y > 10'd364) &&(y <10'd381) )||
    ( (x==  10'd469) &&(y > 10'd364) &&(y <10'd391) )||
    ( (x==  10'd469) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x==  10'd470) &&(y > 10'd361) &&(y <10'd399) )||
    ( (x==  10'd470) &&(y > 10'd349) &&(y <10'd392) )||
    ( (x==  10'd471) &&(y > 10'd321) &&(y <10'd380) )||
    ( (x== 10'd471) &&(y > 10'd397) &&(y <10'd399) )||
    ( (x==  10'd472) &&(y > 10'd321) &&(y <10'd323) )||
    ( (x==  10'd472) &&(y > 10'd325) &&(y <10'd377) )||
    ( (x==  10'd473) &&(y > 10'd321) &&(y <10'd323) )||
    ( (x==  10'd473) &&(y > 10'd325) &&(y <10'd377) )||
    ( (x==  10'd474) &&(y > 10'd321) &&(y <10'd374) )||
    ( (x==  10'd475) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd475) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd475) &&(y > 10'd354) &&(y <10'd357) )||
    ( (x==  10'd476) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd476) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd476) &&(y > 10'd354) &&(y <10'd357) )||
    ( (x==  10'd477) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd477) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x== 10'd477) &&(y > 10'd354) &&(y <10'd360) )||
    ( (x==   10'd478) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd478) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x== 10'd478) &&(y > 10'd355) &&(y <10'd360) )||
    ( (x==  10'd479) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd479) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==   10'd480) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd480) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd481) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==   10'd481) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==   10'd482) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==   10'd482) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==   10'd483) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd483) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd484) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==   10'd484) &&(y > 10'd347) &&(y <10'd350) )||
    ( (x==  10'd485) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd486) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==  10'd487) &&(y > 10'd321) &&(y <10'd347) )||
    ( (x==   10'd488) &&(y > 10'd324) &&(y <10'd347) )||
    ( (x==   10'd489) &&(y > 10'd324) &&(y <10'd347) )||
    ( (x==   10'd490) &&(y > 10'd324) &&(y <10'd347) ) ||
    ( (x== 10'd582) &&(y > 10'd415) &&(y <10'd435) )|| //dino5
    ( (x== 10'd583) &&(y > 10'd418) &&(y <10'd438) )||
    ( (x== 10'd584) &&(y > 10'd421) &&(y <10'd441 ))||
    ( (x== 10'd585) &&(y > 10'd424) &&(y <10'd441 ))||
    ( (x== 10'd586) &&(y > 10'd424) &&(y <10'd441 ))||
    ( (x== 10'd587) &&(y > 10'd424) &&(y <10'd451 ))||
    ( (x== 10'd588) &&(y > 10'd421) &&(y <10'd459 ))||
    ( (x== 10'd589) &&(y > 10'd418) &&(y <10'd455 ))||
    ( (x== 10'd589) &&(y > 10'd457) &&(y <10'd459 ))||
    ( (x== 10'd590) &&(y > 10'd415) &&(y <10'd452) )||
    ( (x== 10'd591) &&(y > 10'd415) &&(y <10'd452) )||
    ( (x== 10'd592) &&(y > 10'd412) &&(y <10'd449) )||
    ( (x==  10'd593) &&(y > 10'd412) &&(y <10'd449) )||
    ( (x==  10'd594) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x==  10'd595) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x== 10'd596) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x== 10'd596) &&(y > 10'd424) &&(y <10'd441) )||
    ( (x==  10'd597) &&(y > 10'd424) &&(y <10'd451) )||
    ( (x==  10'd597) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x==  10'd598) &&(y > 10'd421) &&(y <10'd459) )||
    ( (x==  10'd598) &&(y > 10'd409) &&(y <10'd452) )||
    ( (x==  10'd599) &&(y > 10'd381) &&(y <10'd440) )||
    ( (x== 10'd599) &&(y > 10'd457) &&(y <10'd459) )||
    ( (x==  10'd600) &&(y > 10'd381) &&(y <10'd383) )||
    ( (x==  10'd600) &&(y > 10'd385) &&(y <10'd437) )||
    ( (x==  10'd601) &&(y > 10'd381) &&(y <10'd383) )||
    ( (x==  10'd601) &&(y > 10'd385) &&(y <10'd437) )||
    ( (x==  10'd602) &&(y > 10'd381) &&(y <10'd434) )||
    ( (x==  10'd603) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd603) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd603) &&(y > 10'd414) &&(y <10'd417) )||
    ( (x==  10'd604) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd604) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd604) &&(y > 10'd414) &&(y <10'd417) )||
    ( (x==  10'd605) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd605) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x== 10'd605) &&(y > 10'd414) &&(y <10'd420) )||
    ( (x==   10'd606) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd606) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x== 10'd606) &&(y > 10'd415) &&(y <10'd420) )||
    ( (x==  10'd607) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd607) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==   10'd608) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd608) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd609) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==   10'd609) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==   10'd610) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==   10'd610) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==   10'd611) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd611) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd612) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==   10'd612) &&(y > 10'd407) &&(y <10'd410) )||
    ( (x==  10'd613) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd614) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==  10'd615) &&(y > 10'd381) &&(y <10'd407) )||
    ( (x==   10'd616) &&(y > 10'd384) &&(y <10'd407) )||
    ( (x==   10'd617) &&(y > 10'd384) &&(y <10'd407) )||
    ( (x==   10'd618) &&(y > 10'd384) &&(y <10'd407) ) ||
    ( (x==   10'd87) &&(y > 10'd40) &&(y <10'd111) ) ||//S_left
    ( (x==   10'd88) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd89) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd90) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd91) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd92) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd93) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd94) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd95) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd96) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd97) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd98) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd99) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd100) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd101) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd102) &&(y > 10'd40) &&(y <10'd111) ) ||
    ( (x==   10'd87) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd88) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd89) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd90) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd91) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd92) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd93) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd94) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd95) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd96) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd97) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd98) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd99) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd100) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd101) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd102) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd103) &&(y > 10'd40) &&(y <10'd56) ) ||//S_middle
    ( (x==   10'd104) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd105) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd106) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd107) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd108) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd109) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd110) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd111) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd112) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd113) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd114) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd115) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd116) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd117) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd118) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd119) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd120) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd121) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd122) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd123) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd124) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd125) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd126) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd127) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd128) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd129) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd130) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd131) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd132) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd133) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd134) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd135) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd136) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd137) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd138) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd139) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd140) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd141) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd142) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd143) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd144) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd145) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd146) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd147) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd103) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd104) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd105) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd106) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd107) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd108) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd109) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd110) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd111) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd112) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd113) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd114) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd115) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd116) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd117) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd118) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd119) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd120) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd121) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd122) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd123) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd124) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd125) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd126) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd127) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd128) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd129) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd130) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd131) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd132) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd133) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd134) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd135) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd136) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd137) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd138) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd139) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd140) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd141) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd142) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd143) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd144) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd145) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd146) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd147) &&(y > 10'd95) &&(y <10'd111) ) ||
    ( (x==   10'd103) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd104) &&(y > 10'd144) &&(y <10'd160 )) ||
    ( (x==   10'd105) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd106) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd107) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd108) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd109) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd110) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd111) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd112) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd113) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd114) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd115) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd116) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd117) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd118) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd119) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd120) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd121) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd122) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd123) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd124) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd125) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd126) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd127) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd128) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd129) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd130) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd131) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd132) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd133) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd134) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd135) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd136) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd137) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd138) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd139) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd140) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd141) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd142) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd143) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd144) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd145) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd146) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd147) &&(y > 10'd144) &&(y <10'd160) ) ||
    ( (x==   10'd148) &&(y > 10'd40) &&(y <10'd56) ) ||//S_right
    ( (x==   10'd149) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd150) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd151) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd152) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd153) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd154) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd155) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd156) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd157) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd158) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd159) &&(y > 10'd40) &&(y <10'd56) ) ||
    ( (x==   10'd148) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd149) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd150) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd151) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd152) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd153) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd154) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd155) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd156) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd157) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd158) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (x==   10'd159) &&(y > 10'd95) &&(y <10'd160) ) ||
    ( (y==   10'd41) &&(x > 10'd195) &&(x <10'd265) ) ||//T_up
    ( (y==   10'd42) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd43) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd44) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd45) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd46) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd47) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd48) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd49) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd50) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd51) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd52) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd53) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd54) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd55) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (y==   10'd56) &&(x > 10'd195) &&(x <10'd265) ) ||
    ( (x==   10'd222) &&(y > 10'd56) &&(y <10'd160) ) ||//T_down
    ( (x==   10'd223) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd224) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd225) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd226) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd227) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd228) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd229) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd230) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd231) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd232) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd233) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd234) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd235) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd236) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd237) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd238) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd280) &&(y > 10'd40) &&(y <10'd160) ) ||//A_left
    ( (x==   10'd281) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd282) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd283) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd284) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd285) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd286) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd287) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd288) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd289) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd290) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd291) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd292) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd293) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd294) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd295) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (y==   10'd41) &&(x > 10'd295) &&(x <10'd345) ) ||//A_middle_up
    ( (y==   10'd42) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd43) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd44) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd45) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd46) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd47) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd48) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd49) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd50) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd51) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd52) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd53) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd54) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd55) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd56) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd101) &&(x > 10'd295) &&(x <10'd345) ) ||//A_middle_middle
    ( (y==   10'd102) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd103) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd104) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd105) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd106) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd107) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd108) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd109) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd110) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd111) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd112) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd113) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd114) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd115) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (y==   10'd116) &&(x > 10'd295) &&(x <10'd345) ) ||
    ( (x==   10'd345) &&(y > 10'd40) &&(y <10'd160) ) ||//A_right
    ( (x==   10'd346) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd347) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd348) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd349) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd350) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd351) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd352) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd353) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd354) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd355) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd356) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd357) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd358) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd359) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd375) &&(y > 10'd40) &&(y <10'd160) ) ||//R_left
    ( (x==   10'd376) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd377) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd378) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd379) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd380) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd381) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd382) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd383) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd384) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd385) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd386) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd387) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd388) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd389) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (x==   10'd390) &&(y > 10'd40) &&(y <10'd160) ) ||
    ( (y==   10'd41) &&(x > 10'd390) &&(x <10'd440) ) ||//R_middle_up
    ( (y==   10'd42) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd43) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd44) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd45) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd46) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd47) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd48) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd49) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd50) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd51) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd52) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd53) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd54) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd55) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd56) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd101) &&(x > 10'd390) &&(x <10'd440) ) ||//R_middle_middle
    ( (y==   10'd102) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd103) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd104) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd105) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd106) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd107) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd108) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd109) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd110) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd111) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd112) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd113) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd114) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd115) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (y==   10'd116) &&(x > 10'd390) &&(x <10'd440) ) ||
    ( (x==   10'd440) &&(y > 10'd40) &&(y <10'd117) ) ||//R_right
    ( (x==   10'd441) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd442) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd443) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd444) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd445) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd446) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd447) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd448) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd449) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd450) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd451) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd452) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd453) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd454) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd455) &&(y > 10'd40) &&(y <10'd117) ) ||
    ( (x==   10'd391) &&(y > 10'd116) &&(y <10'd134) ) ||//R_slash
    ( (x==   10'd392) &&(y > 10'd116) &&(y <10'd134) ) ||
    ( (x==   10'd393) &&(y > 10'd116) &&(y <10'd134) )||
    ( (x==   10'd394) &&(y > 10'd116) &&(y <10'd135) )||
    ( (x==   10'd395) &&(y > 10'd116) &&(y <10'd135) )||
    ( (x==   10'd396) &&(y > 10'd116) &&(y <10'd136) )||
    ( (x==   10'd397) &&(y > 10'd117) &&(y <10'd137) )||
    ( (x==   10'd398) &&(y > 10'd117) &&(y <10'd137) )||
    ( (x==   10'd399) &&(y > 10'd117) &&(y <10'd137) )||
    ( (x==   10'd400) &&(y > 10'd118) &&(y <10'd138) )||
    ( (x==   10'd401) &&(y > 10'd118) &&(y <10'd138) )||
    ( (x==   10'd402) &&(y > 10'd119) &&(y <10'd139) )||
    ( (x==   10'd403) &&(y > 10'd119) &&(y <10'd139) )||
    ( (x==   10'd404) &&(y > 10'd119) &&(y <10'd139) )||
    ( (x==   10'd405) &&(y > 10'd120) &&(y <10'd140) )||
    ( (x==   10'd406) &&(y > 10'd120) &&(y <10'd140) )||
    ( (x==   10'd407) &&(y > 10'd121) &&(y <10'd141) )||
    ( (x==   10'd408) &&(y > 10'd121) &&(y <10'd141) )||
    ( (x==   10'd409) &&(y > 10'd121) &&(y <10'd141) )||
    ( (x==   10'd410) &&(y > 10'd122) &&(y <10'd142) )||
    ( (x==   10'd411) &&(y > 10'd122) &&(y <10'd142) )||
    ( (x==   10'd412) &&(y > 10'd123) &&(y <10'd143) )||
    ( (x==   10'd413) &&(y > 10'd123) &&(y <10'd143) )||
    ( (x==   10'd414) &&(y > 10'd123) &&(y <10'd143) )||
    ( (x==   10'd415) &&(y > 10'd124) &&(y <10'd144) )||
    ( (x==   10'd416) &&(y > 10'd124) &&(y <10'd144) )||
    ( (x==   10'd417) &&(y > 10'd125) &&(y <10'd145) )||
    ( (x==   10'd418) &&(y > 10'd125) &&(y <10'd145) )||
    ( (x==   10'd419) &&(y > 10'd125) &&(y <10'd145) )||
    ( (x==   10'd420) &&(y > 10'd126) &&(y <10'd146) ) ||
    ( (x==   10'd421) &&(y > 10'd126) &&(y <10'd146) ) ||
    ( (x==   10'd422) &&(y > 10'd127) &&(y <10'd147) )||
    ( (x==   10'd423) &&(y > 10'd127) &&(y <10'd147) )||
    ( (x==   10'd424) &&(y > 10'd127) &&(y <10'd147) )||
    ( (x==   10'd425) &&(y > 10'd128) &&(y <10'd148) )||
    ( (x==   10'd426) &&(y > 10'd128) &&(y <10'd148) )||
    ( (x==   10'd427) &&(y > 10'd129) &&(y <10'd149) )||
    ( (x==   10'd428) &&(y > 10'd129) &&(y <10'd149) )||
    ( (x==   10'd429) &&(y > 10'd129) &&(y <10'd149) )||
    ( (x==   10'd430) &&(y > 10'd130) &&(y <10'd150) )||
    ( (x==   10'd431) &&(y > 10'd130) &&(y <10'd150) )||
    ( (x==   10'd432) &&(y > 10'd131) &&(y <10'd151) )||
    ( (x==   10'd433) &&(y > 10'd131) &&(y <10'd151) )||
     ( (x==   10'd434) &&(y > 10'd131) &&(y <10'd151) )||
    ( (x==   10'd435) &&(y > 10'd132) &&(y <10'd152) )||
    ( (x==   10'd436) &&(y > 10'd132) &&(y <10'd152) )||
    ( (x==   10'd437) &&(y > 10'd133) &&(y <10'd153) ) ||
    ( (x==   10'd438) &&(y > 10'd133) &&(y <10'd153) ) ||
    ( (x==   10'd439) &&(y > 10'd133) &&(y <10'd153) ) ||
    ( (x==   10'd440) &&(y > 10'd134) &&(y <10'd154) )||
    ( (x==   10'd441) &&(y > 10'd134) &&(y <10'd154) )||
    ( (x==   10'd442) &&(y > 10'd135) &&(y <10'd155) )||
    ( (x==   10'd443) &&(y > 10'd135) &&(y <10'd155) )||
    ( (x==   10'd444) &&(y > 10'd135) &&(y <10'd155) )||
    ( (x==   10'd445) &&(y > 10'd136) &&(y <10'd156) )||
    ( (x==   10'd446) &&(y > 10'd136) &&(y <10'd156) )||
    ( (x==   10'd447) &&(y > 10'd137) &&(y <10'd157) )||
    ( (x==   10'd448) &&(y > 10'd137) &&(y <10'd157) )||
    ( (x==   10'd449) &&(y > 10'd137) &&(y <10'd157) )||
    ( (x==   10'd450) &&(y > 10'd138) &&(y <10'd158) )||
    ( (x==   10'd451) &&(y > 10'd138) &&(y <10'd158) )||
    ( (x==   10'd452) &&(y > 10'd139) &&(y <10'd159) )||
    ( (x==   10'd453) &&(y > 10'd139) &&(y <10'd159) )||
    ( (x==   10'd454) &&(y > 10'd139) &&(y <10'd159) )||
    ( (x==   10'd455) &&(y > 10'd140) &&(y <10'd160) ) ||
    ( (x==   10'd456) &&(y > 10'd140) &&(y <10'd160) ) ||
    ( (y==   10'd41) &&(x > 10'd483) &&(x <10'd553) ) ||//T2_up
    ( (y==   10'd42) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd43) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd44) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd45) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd46) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd47) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd48) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd49) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd50) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd51) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd52) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd53) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd54) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd55) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (y==   10'd56) &&(x > 10'd483) &&(x <10'd553) ) ||
    ( (x==   10'd510) &&(y > 10'd56) &&(y <10'd160) ) ||//T2_down
    ( (x==   10'd511) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd512) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd513) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd514) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd515) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd516) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd517) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd518) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd519) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd520) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd521) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd522) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd523) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd524) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd525) &&(y > 10'd56) &&(y <10'd160) ) ||
    ( (x==   10'd526) &&(y > 10'd56) &&(y <10'd160) ) 
     
    ;
    
    assign bird_draw =  
    ( (x== (bird_x + 10'd1)) &&(y > (bird_y+10'd17)) &&(y <bird_y+10'd20) )||//head
    ( (x== (bird_x + 10'd2)) &&(y > (bird_y+10'd17)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd3)) &&(y > (bird_y+10'd15)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd4)) &&(y > (bird_y+10'd15)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd5)) &&(y > (bird_y+10'd13)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd6)) &&(y > (bird_y+10'd13)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd7)) &&(y > (bird_y+10'd11)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd8)) &&(y > (bird_y+10'd11)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd9)) &&(y > (bird_y+10'd7)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd10)) &&(y > (bird_y+10'd7)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd11)) &&(y > (bird_y+10'd7)) &&(y <bird_y+10'd20) )||
    ( (x== (bird_x + 10'd12)) &&(y > (bird_y+10'd13)) &&(y <bird_y+10'd22) )||//neck
    ( (x== (bird_x + 10'd13)) &&(y > (bird_y+10'd1)) &&(y <bird_y+10'd8) )||
    ( (x== (bird_x + 10'd13)) &&(y > (bird_y+10'd15)) &&(y <bird_y+10'd24) )||
    ( (x== (bird_x + 10'd14)) &&(y > (bird_y+10'd5)) &&(y <bird_y+10'd26) )||//body
    ( (x== (bird_x + 10'd15)) &&(y > (bird_y+10'd5)) &&(y <bird_y+10'd26) )||
    ( (x== (bird_x + 10'd16)) &&(y > (bird_y+10'd7)) &&(y <bird_y+10'd28) )||
    ( (x== (bird_x + 10'd17)) &&(y > (bird_y+10'd7)) &&(y <bird_y+10'd28) )||
    ( (x== (bird_x + 10'd18)) &&(y > (bird_y+10'd9)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd19)) &&(y > (bird_y+10'd9)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd20)) &&(y > (bird_y+10'd11)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd21)) &&(y > (bird_y+10'd11)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd22)) &&(y > (bird_y+10'd13)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd23)) &&(y > (bird_y+10'd13)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd24)) &&(y > (bird_y+10'd15)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd25)) &&(y > (bird_y+10'd15)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd26)) &&(y > (bird_y+10'd17)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd27)) &&(y > (bird_y+10'd17)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd28)) &&(y > (bird_y+10'd19)) &&(y <bird_y+10'd30) )||
    ( (x== (bird_x + 10'd28)) &&(y > (bird_y+10'd19)) &&(y <bird_y+10'd30) ) ||
    ( (x== (bird_x + 10'd29)) &&(y > (bird_y+10'd23)) &&(y <bird_y+10'd27) ) ||//tail
    ( (x== (bird_x + 10'd30)) &&(y > (bird_y+10'd23)) &&(y <bird_y+10'd27) ) ||
    ( (x== (bird_x + 10'd31)) &&(y > (bird_y+10'd23)) &&(y <bird_y+10'd26) ) ||
    ( (x== (bird_x + 10'd31)) &&(y > (bird_y+10'd26)) &&(y <bird_y+10'd29) ) ||
    ( (x== (bird_x + 10'd32)) &&(y > (bird_y+10'd23)) &&(y <bird_y+10'd26) ) ||
    ( (x== (bird_x + 10'd32)) &&(y > (bird_y+10'd26)) &&(y <bird_y+10'd29) ) ||
    ( (x== (bird_x + 10'd33)) &&(y > (bird_y+10'd23)) &&(y <bird_y+10'd26) ) ||
    ( (x== (bird_x + 10'd34)) &&(y > (bird_y+10'd23)) &&(y <bird_y+10'd26) ) 
    ;

    always @(posedge clk)begin
        if(rst)
             pixel <= 12'hfff;
        else begin
            if(state == 2'b00)begin//start == stop
                if(black)
                pixel <= 12'h000;
                else
                pixel <= 12'hfff;
            end else if(state == 2'b01)begin//game
                if( obtacle_draw )
                    pixel <= 12'h000;
                else if(dino_draw)
                    pixel <= 12'h000;
                else if(bird_draw)
                    pixel <= 12'h000;
                else begin
                    if(sun)
                        pixel <= 12'hfa0;
                    else if(cloud)
                        pixel <= 12'hfff;
                    else if(y <= 180)
                        pixel <= 12'h0ff;
                    else
                        pixel <= 12'hfff;
                end
            end else begin
                pixel <= 12'h000;
            end
            
        end
    end
 
           
endmodule
